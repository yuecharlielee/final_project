`include "global.v"

module mem_addr_gen(
    h_cnt, v_cnt,
    x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9, 
    y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7, y_8, y_9, 
    s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9,
    pixel_addr
    );
    
    input [9:0] h_cnt;
    input [9:0] v_cnt;

    input [9:0] x_0, x_1, x_2, x_3, x_4, x_5, x_6, x_7, x_8, x_9;
    input [9:0] y_0, y_1, y_2, y_3, y_4, y_5, y_6, y_7, y_8, y_9;
    input [9:0] s_0, s_1, s_2, s_3, s_4, s_5, s_6, s_7, s_8, s_9;

    output reg [16:0] pixel_addr;

     
    wire [19:0] h_cnt_rs;
    wire [19:0] v_cnt_rs;

    assign h_cnt_rs = h_cnt >> 1; 
    assign v_cnt_rs = v_cnt >> 1; 

    wire in_circle_0 = (h_cnt_rs - x_0) * (h_cnt_rs - x_0) + (v_cnt_rs - y_0) * (v_cnt_rs - y_0) < `ball_size_0 * `ball_size_0;
    wire in_circle_1 = (h_cnt_rs - x_1) * (h_cnt_rs - x_1) + (v_cnt_rs - y_1) * (v_cnt_rs - y_1) < `ball_size_0 * `ball_size_0;
    wire in_circle_2 = (h_cnt_rs - x_2) * (h_cnt_rs - x_2) + (v_cnt_rs - y_2) * (v_cnt_rs - y_2) < `ball_size_0 * `ball_size_0;
    wire in_circle_3 = (h_cnt_rs - x_3) * (h_cnt_rs - x_3) + (v_cnt_rs - y_3) * (v_cnt_rs - y_3) < `ball_size_0 * `ball_size_0;
    wire in_circle_4 = (h_cnt_rs - x_4) * (h_cnt_rs - x_4) + (v_cnt_rs - y_4) * (v_cnt_rs - y_4) < `ball_size_0 * `ball_size_0;
    wire in_circle_5 = (h_cnt_rs - x_5) * (h_cnt_rs - x_5) + (v_cnt_rs - y_5) * (v_cnt_rs - y_5) < `ball_size_0 * `ball_size_0;
    wire in_circle_6 = (h_cnt_rs - x_6) * (h_cnt_rs - x_6) + (v_cnt_rs - y_6) * (v_cnt_rs - y_6) < `ball_size_0 * `ball_size_0;
    wire in_circle_7 = (h_cnt_rs - x_7) * (h_cnt_rs - x_7) + (v_cnt_rs - y_7) * (v_cnt_rs - y_7) < `ball_size_0 * `ball_size_0;
    wire in_circle_8 = (h_cnt_rs - x_8) * (h_cnt_rs - x_8) + (v_cnt_rs - y_8) * (v_cnt_rs - y_8) < `ball_size_0 * `ball_size_0;
    wire in_circle_9 = (h_cnt_rs - x_9) * (h_cnt_rs - x_9) + (v_cnt_rs - y_9) * (v_cnt_rs - y_9) < `ball_size_0 * `ball_size_0;
    //wire in_circle_2 = (h_cnt_rs - x_2) * (h_cnt_rs - x_2) + (v_cnt_rs - y_2) * (v_cnt_rs - y_2) < size_2 * size_2;

    wire in_circle = in_circle_0 || in_circle_1 || in_circle_2 || in_circle_3 || in_circle_4 || in_circle_5 || in_circle_6 || in_circle_7 || in_circle_8 || in_circle_9; 

    always @ (*) begin
        if(in_circle) begin
            pixel_addr = 17'd4000;
        end
        else begin
            if(v_cnt_rs <= `up_bound || h_cnt_rs <= `left_bound || h_cnt_rs >= `right_bound) begin
                pixel_addr = 0;
            end
            else begin
                pixel_addr = ((h_cnt_rs)+320*(v_cnt_rs))% 76800;
            end
        end
        
    end
    
    always @(*) begin
        
    end
    
endmodule
